library verilog;
use verilog.vl_types.all;
entity eight_one_mux_tb is
end eight_one_mux_tb;
